* Spice description of cronometro_cougar
* Spice driver version -1218054087
* Date ( dd/mm/yyyy hh:mm:ss ): 22/04/2018 at  2:20:08

* INTERF ctrl dmin[0] dmin[1] dmin[2] dseg[0] dseg[1] dseg[2] rlj rst 
* INTERF umin[0] umin[1] umin[2] umin[3] useg[0] useg[1] useg[2] useg[3] vdd 
* INTERF vss 


.subckt cronometro_cougar 133 530 525 524 149 187 185 515 488 521 506 503 492 
+ 27 22 25 20 534 487 
* NET 11 = memuseg_3_ins.sff_s
* NET 13 = memuseg_3_ins.y
* NET 14 = memuseg_3_ins.sff_m
* NET 17 = memuseg_3_ins.u
* NET 18 = memuseg_3_ins.ckr
* NET 19 = memuseg_3_ins.nckr
* NET 20 = useg[3]
* NET 22 = useg[1]
* NET 25 = useg[2]
* NET 26 = aux19
* NET 27 = useg[0]
* NET 29 = no2_x1_9_sig
* NET 30 = no2_x1_10_sig
* NET 36 = maquina_0_ins.sff_m
* NET 37 = maquina_0_ins.sff_s
* NET 38 = maquina_0_ins.y
* NET 39 = oa2a22_x2_4_sig
* NET 41 = maquina_0_ins.u
* NET 42 = maquina_0_ins.ckr
* NET 43 = maquina_0_ins.nckr
* NET 57 = a3_x2_3_sig
* NET 58 = oa22_x2_4_sig
* NET 60 = oa22_x2_5_sig
* NET 69 = nao22_x1_4_sig
* NET 72 = nao22_x1_5_sig
* NET 74 = a2_x2_6_sig
* NET 82 = not_aux21
* NET 86 = not_aux18
* NET 89 = not_maquina[0]
* NET 90 = no2_x1_7_sig
* NET 91 = maquina[0]
* NET 92 = no2_x1_8_sig
* NET 96 = maquina[1]
* NET 99 = maquina_1_ins.y
* NET 101 = maquina_1_ins.sff_m
* NET 102 = maquina_1_ins.sff_s
* NET 104 = oa2a22_x2_3_sig
* NET 105 = maquina_1_ins.u
* NET 107 = maquina_1_ins.nckr
* NET 108 = maquina_1_ins.ckr
* NET 112 = no3_x1_5_sig
* NET 113 = aux23
* NET 114 = a3_x2_2_sig
* NET 118 = mbk_buf_not_aux0
* NET 121 = memuseg_1_ins.y
* NET 122 = memuseg_1_ins.sff_m
* NET 124 = memuseg_1_ins.sff_s
* NET 125 = oa22_x2_3_sig
* NET 126 = memuseg_1_ins.u
* NET 128 = memuseg_1_ins.ckr
* NET 129 = memuseg_1_ins.nckr
* NET 130 = aux24
* NET 133 = ctrl
* NET 134 = not_ctrl
* NET 135 = not_aux20
* NET 136 = not_aux22
* NET 139 = memuseg_0_ins.y
* NET 140 = memuseg_0_ins.sff_s
* NET 141 = memuseg_0_ins.sff_m
* NET 143 = nao22_x1_3_sig
* NET 144 = memuseg_0_ins.nckr
* NET 145 = memuseg_0_ins.u
* NET 147 = memuseg_0_ins.ckr
* NET 149 = dseg[0]
* NET 157 = na2_x1_sig
* NET 158 = not_aux23
* NET 162 = not_aux19
* NET 166 = o3_x2_4_sig
* NET 167 = o3_x2_3_sig
* NET 168 = na2_x1_2_sig
* NET 171 = memuseg[2]
* NET 173 = memuseg_2_ins.y
* NET 175 = memuseg_2_ins.sff_s
* NET 177 = na3_x1_sig
* NET 178 = memuseg_2_ins.ckr
* NET 179 = memuseg_2_ins.u
* NET 180 = memuseg_2_ins.sff_m
* NET 182 = memuseg[0]
* NET 183 = memuseg_2_ins.nckr
* NET 185 = dseg[2]
* NET 187 = dseg[1]
* NET 191 = inv_x2_2_sig
* NET 192 = not_memuseg[1]
* NET 197 = no3_x1_4_sig
* NET 201 = memuseg[3]
* NET 202 = no2_x1_5_sig
* NET 203 = not_aux0
* NET 204 = mbk_buf_memuseg[2]
* NET 205 = memuseg[1]
* NET 206 = not_memuseg[3]
* NET 210 = mbk_buf_not_memuseg[2]
* NET 211 = not_memuseg[2]
* NET 216 = memdseg_2_ins.ckr
* NET 217 = memdseg_2_ins.u
* NET 219 = memdseg_2_ins.nckr
* NET 220 = oa2a22_x2_2_sig
* NET 232 = mx2_x2_sig
* NET 233 = memdseg_1_ins.u
* NET 234 = memdseg_1_ins.ckr
* NET 235 = memdseg_1_ins.nckr
* NET 245 = memdseg_2_ins.sff_s
* NET 246 = memdseg_2_ins.y
* NET 247 = memdseg_2_ins.sff_m
* NET 257 = memdseg_1_ins.sff_s
* NET 258 = memdseg_1_ins.y
* NET 259 = memdseg_1_ins.sff_m
* NET 264 = memdseg_0_ins.sff_s
* NET 265 = memdseg_0_ins.y
* NET 267 = memdseg_0_ins.u
* NET 269 = memdseg_0_ins.sff_m
* NET 270 = memdseg_0_ins.ckr
* NET 271 = a3_x2_sig
* NET 272 = oa22_x2_2_sig
* NET 273 = memdseg_0_ins.nckr
* NET 274 = no4_x1_sig
* NET 277 = not_memuseg[0]
* NET 278 = no3_x1_sig
* NET 281 = not_aux8
* NET 282 = inv_x2_sig
* NET 285 = memumin_0_ins.sff_s
* NET 286 = memumin_0_ins.y
* NET 289 = memumin_0_ins.ckr
* NET 290 = memumin_0_ins.u
* NET 291 = memumin_0_ins.sff_m
* NET 292 = memumin_0_ins.nckr
* NET 294 = aux30
* NET 297 = oa2ao222_x2_3_sig
* NET 299 = memdseg[2]
* NET 300 = a2_x2_5_sig
* NET 303 = not_memdseg[2]
* NET 304 = a2_x2_4_sig
* NET 307 = memdseg[1]
* NET 309 = nxr2_x1_2_sig
* NET 312 = no2_x1_6_sig
* NET 325 = aux28
* NET 337 = mbk_buf_not_aux2
* NET 339 = memdseg[0]
* NET 340 = not_aux2
* NET 343 = mbk_buf_aux3
* NET 345 = memdmin_0_ins.sff_s
* NET 346 = aux3
* NET 347 = memdmin_0_ins.sff_m
* NET 348 = memdmin_0_ins.ckr
* NET 350 = memdmin_0_ins.y
* NET 354 = memdmin_0_ins.nckr
* NET 355 = memdmin_0_ins.u
* NET 363 = oa2a22_x2_sig
* NET 365 = xr2_x1_sig
* NET 369 = aux27
* NET 371 = a2_x2_sig
* NET 377 = memdmin_1_ins.sff_s
* NET 379 = memdmin_1_ins.sff_m
* NET 380 = memdmin_1_ins.ckr
* NET 382 = memdmin_1_ins.y
* NET 384 = memdmin_1_ins.u
* NET 385 = oa2ao222_x2_sig
* NET 386 = memdmin_1_ins.nckr
* NET 389 = nao22_x1_2_sig
* NET 393 = o3_x2_2_sig
* NET 396 = not_aux3
* NET 398 = memumin_3_ins.sff_s
* NET 400 = oa22_x2_sig
* NET 401 = memumin_3_ins.y
* NET 402 = memumin_3_ins.sff_m
* NET 405 = memumin_3_ins.nckr
* NET 406 = memumin_3_ins.ckr
* NET 407 = memumin_3_ins.u
* NET 409 = not_aux6
* NET 412 = a2_x2_3_sig
* NET 413 = aux25
* NET 414 = aux26
* NET 419 = memdmin_2_ins.sff_s
* NET 420 = memdmin_2_ins.y
* NET 422 = memdmin_2_ins.sff_m
* NET 423 = oa2ao222_x2_2_sig
* NET 424 = memdmin_2_ins.u
* NET 426 = memdmin_2_ins.ckr
* NET 427 = memdmin_2_ins.nckr
* NET 446 = not_aux17
* NET 447 = not_memumin[3]
* NET 448 = nao2o22_x1_sig
* NET 451 = not_memumin[2]
* NET 454 = no2_x1_2_sig
* NET 456 = not_aux16
* NET 457 = o3_x2_sig
* NET 459 = not_memumin[1]
* NET 461 = memumin_1_ins.sff_s
* NET 463 = memumin_1_ins.y
* NET 464 = memumin_1_ins.sff_m
* NET 469 = nao22_x1_sig
* NET 470 = memumin_1_ins.nckr
* NET 471 = memumin_1_ins.u
* NET 472 = memumin_1_ins.ckr
* NET 477 = mbk_buf_not_aux8
* NET 478 = nxr2_x1_sig
* NET 479 = no3_x1_3_sig
* NET 480 = aux8
* NET 481 = ao22_x2_sig
* NET 484 = no3_x1_2_sig
* NET 486 = no2_x1_sig
* NET 487 = vss
* NET 488 = rst
* NET 489 = memumin[3]
* NET 490 = not_aux29
* NET 492 = umin[3]
* NET 493 = inv_x2_3_sig
* NET 494 = not_rst
* NET 495 = no2_x1_4_sig
* NET 499 = not_aux14
* NET 500 = no2_x1_3_sig
* NET 503 = umin[2]
* NET 504 = memumin[1]
* NET 506 = umin[1]
* NET 508 = memumin[2]
* NET 510 = memumin_2_ins.sff_s
* NET 511 = memumin_2_ins.y
* NET 513 = memumin_2_ins.sff_m
* NET 514 = oa2ao222_x2_4_sig
* NET 515 = rlj
* NET 516 = memumin_2_ins.nckr
* NET 517 = memumin_2_ins.u
* NET 518 = memumin_2_ins.ckr
* NET 519 = memumin[0]
* NET 521 = umin[0]
* NET 522 = memdmin[2]
* NET 524 = dmin[2]
* NET 525 = dmin[1]
* NET 527 = a2_x2_2_sig
* NET 528 = memdmin[1]
* NET 530 = dmin[0]
* NET 531 = memdmin[0]
* NET 532 = not_memdmin[0]
* NET 534 = vdd
Mtr_01058 525 526 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01057 534 528 526 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01056 527 529 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01055 534 532 529 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01054 529 528 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01053 521 520 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01052 534 519 520 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01051 530 533 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01050 534 531 533 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01049 532 531 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01048 493 490 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01047 492 491 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01046 534 489 491 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01045 507 508 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01044 510 518 507 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01043 511 516 510 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01042 513 516 512 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01041 512 511 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01040 509 518 513 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01039 516 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01038 534 516 518 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01037 517 514 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01036 534 517 509 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01035 534 510 508 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01034 508 510 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01033 511 513 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01032 506 505 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01031 534 504 505 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01030 524 523 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01029 534 522 523 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01028 501 508 500 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01027 534 499 501 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01026 503 502 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01025 534 508 502 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_01024 514 497 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01023 496 500 498 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01022 496 494 534 534 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_01021 534 493 496 534 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_01020 498 495 497 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01019 497 504 496 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01018 494 488 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_01017 534 477 441 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01016 440 478 479 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01015 441 486 440 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01014 445 532 486 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01013 534 528 445 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01012 534 482 481 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01011 482 480 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01010 534 484 442 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01009 442 527 482 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01008 534 522 443 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01007 444 532 484 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01006 443 528 444 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01005 534 474 439 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01004 439 476 478 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01003 439 531 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01002 478 522 439 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_01001 534 531 476 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_01000 474 522 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00999 534 504 434 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00998 434 499 433 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00997 433 454 455 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00996 457 455 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00995 534 457 469 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00994 435 456 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00993 469 459 435 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00992 436 504 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00991 461 472 436 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00990 463 470 461 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00989 464 470 438 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00988 438 463 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00987 437 472 464 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00986 470 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00985 534 470 472 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00984 471 469 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00983 534 471 437 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00982 534 461 504 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00981 504 461 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00980 463 464 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00979 428 447 454 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00978 534 508 428 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00977 431 451 450 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00976 534 504 431 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00975 490 450 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00974 432 456 495 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00973 534 451 432 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00972 448 456 430 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00971 430 447 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00970 429 446 448 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00969 534 490 429 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00968 447 489 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00967 459 504 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00966 418 522 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00965 419 426 418 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00964 420 427 419 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00963 422 427 421 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00962 421 420 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00961 425 426 422 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00960 427 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00959 534 427 426 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00958 424 423 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00957 534 424 425 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00956 534 419 522 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00955 522 419 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00954 420 422 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00953 412 411 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00952 534 522 411 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00951 411 477 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00950 423 417 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00949 415 412 416 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00948 415 413 534 534 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00947 534 522 415 534 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00946 416 479 417 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00945 417 414 415 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00944 409 397 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00943 397 396 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00942 534 489 397 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00941 397 451 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00940 534 459 397 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00939 410 409 413 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00938 534 488 410 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00937 414 408 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00936 534 409 408 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00935 408 494 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00934 451 508 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00933 534 390 400 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00932 391 448 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00931 391 389 390 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00930 390 504 391 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00929 534 489 394 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00928 394 499 395 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00927 395 451 392 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00926 393 392 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00925 399 489 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00924 398 406 399 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00923 401 405 398 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00922 402 405 404 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00921 404 401 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00920 403 406 402 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00919 405 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00918 534 405 406 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00917 407 400 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00916 534 407 403 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00915 534 398 489 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00914 489 398 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00913 401 402 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00912 446 494 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00911 534 489 446 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00910 534 393 389 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00909 388 508 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00908 389 446 388 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00907 371 370 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00906 534 528 370 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00905 370 477 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00904 330 528 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00903 377 380 330 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00902 382 386 377 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00901 379 386 332 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00900 332 382 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00899 333 380 379 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00898 386 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00897 534 386 380 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00896 384 385 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00895 534 384 333 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00894 534 377 528 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00893 528 377 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00892 382 379 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00891 323 365 362 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00890 323 413 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00889 534 531 323 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00888 362 414 323 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00887 363 362 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00886 316 531 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00885 345 348 316 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00884 350 354 345 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00883 347 354 315 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00882 315 350 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00881 318 348 347 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00880 354 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00879 534 354 348 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00878 355 363 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00877 534 355 318 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00876 534 345 531 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00875 531 345 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00874 350 347 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00873 385 373 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00872 329 371 326 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00871 329 413 534 534 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00870 534 528 329 534 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00869 326 481 373 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00868 373 414 329 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00867 534 494 456 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00866 314 477 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00865 456 343 314 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00864 369 367 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00863 534 494 367 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00862 367 396 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00861 358 531 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00860 534 480 357 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00859 365 358 320 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00858 320 480 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00857 320 357 365 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00856 534 531 320 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00855 396 346 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00854 337 335 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00853 534 340 335 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00852 311 337 312 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00851 534 488 311 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00850 324 396 325 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00849 534 488 324 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00848 343 338 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00847 534 346 338 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00846 346 339 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00845 534 340 346 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00844 284 519 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00843 285 289 284 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00842 286 292 285 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00841 291 292 287 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00840 287 286 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00839 288 289 291 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00838 292 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00837 534 292 289 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00836 290 297 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00835 534 290 288 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00834 534 285 519 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00833 519 285 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00832 286 291 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00831 297 296 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00830 302 304 298 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00829 302 325 534 534 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00828 534 519 302 534 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00827 298 300 296 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00826 296 369 302 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00825 534 306 310 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00824 310 308 309 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00823 310 519 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00822 309 307 310 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00821 534 519 308 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00820 306 307 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00819 304 305 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00818 534 303 305 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00817 305 519 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00816 293 369 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00815 534 293 295 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00814 295 299 294 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00813 534 488 280 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00812 279 277 278 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00811 280 282 279 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00810 477 283 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00809 534 281 283 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00808 499 278 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00807 534 274 499 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00806 300 301 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00805 534 299 301 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00804 301 309 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00803 282 339 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00802 263 339 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00801 264 270 263 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00800 265 273 264 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00799 269 273 266 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00798 266 265 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00797 268 270 269 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00796 273 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00795 534 273 270 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00794 267 272 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00793 534 267 268 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00792 534 264 339 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00791 339 264 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00790 265 269 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00789 534 275 272 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00788 276 271 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00787 276 339 275 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00786 275 312 276 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00785 281 480 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00784 188 307 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00783 257 234 188 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00782 258 235 257 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00781 259 235 230 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00780 230 258 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00779 229 234 259 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00778 235 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00777 534 235 234 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00776 233 232 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00775 534 233 229 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00774 534 257 307 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00773 307 257 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00772 258 259 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00771 534 252 232 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00770 224 325 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00769 254 307 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00768 225 307 252 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00767 252 254 224 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00766 534 294 225 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00765 223 307 251 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00764 223 325 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00763 534 299 223 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00762 251 294 223 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00761 220 251 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00760 172 299 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00759 245 216 172 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00758 246 219 245 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00757 247 219 212 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00756 212 246 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00755 215 216 247 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00754 219 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00753 534 219 216 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00752 217 220 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00751 534 217 215 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00750 534 245 299 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00749 299 245 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00748 246 247 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00747 534 339 196 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00746 195 277 197 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00745 196 488 195 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00744 534 197 240 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00743 271 240 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00742 534 210 240 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00741 240 202 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00740 534 281 207 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00739 208 205 209 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00738 209 206 274 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00737 207 204 208 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00736 210 244 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00735 534 211 244 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00734 192 205 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00733 534 203 237 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00732 340 237 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00731 534 201 237 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00730 237 192 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00729 206 201 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00728 198 206 202 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00727 534 205 198 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00726 534 303 190 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00725 189 307 480 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00724 190 191 189 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00723 203 170 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00722 534 211 170 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00721 170 182 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00720 185 184 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00719 534 299 184 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00718 303 299 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00717 187 186 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00716 534 307 186 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00715 191 519 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00714 277 182 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00713 204 169 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00712 534 171 169 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00711 534 162 164 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00710 164 205 163 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00709 163 210 165 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00708 167 165 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00707 534 166 177 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00706 177 167 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00705 177 168 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00704 176 171 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00703 175 178 176 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00702 173 183 175 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00701 180 183 174 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00700 174 173 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00699 181 178 180 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00698 183 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00697 534 183 178 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00696 179 177 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00695 534 179 181 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00694 534 175 171 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00693 171 175 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00692 173 180 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00691 157 201 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00690 534 210 157 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00689 534 158 161 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00688 161 204 159 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00687 159 192 160 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00686 166 160 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00685 534 171 211 534 tp L=1U W=14U AS=28P AD=28P PS=32U PD=32U 
Mtr_00684 211 171 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00683 118 119 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00682 534 203 119 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00681 95 182 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00680 140 147 95 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00679 139 144 140 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00678 141 144 98 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00677 98 139 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00676 103 147 141 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00675 144 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00674 534 144 147 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00673 145 143 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00672 534 145 103 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00671 534 140 182 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00670 182 140 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00669 139 141 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00668 149 148 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00667 534 339 148 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00666 134 133 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00665 67 277 113 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00664 534 162 67 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00663 85 182 132 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00662 534 162 85 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00661 135 132 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00660 130 135 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00659 534 136 130 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00658 534 135 143 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00657 88 136 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00656 143 277 88 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00655 168 130 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00654 534 204 168 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00653 75 205 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00652 124 128 75 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00651 121 129 124 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00650 122 129 78 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00649 78 121 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00648 80 128 122 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00647 129 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00646 534 129 128 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00645 126 125 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00644 534 126 80 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00643 534 124 205 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00642 205 124 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00641 121 122 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00640 534 113 110 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00639 114 110 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00638 534 192 110 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00637 110 157 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00636 158 113 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00635 534 201 64 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00634 63 210 112 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00633 64 158 63 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00632 534 115 125 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00631 70 114 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00630 70 205 115 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00629 115 130 70 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00628 94 89 93 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00627 94 90 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00626 534 91 94 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00625 93 92 94 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00624 104 93 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00623 97 96 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00622 102 108 97 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00621 99 107 102 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00620 101 107 100 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00619 100 99 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00618 106 108 101 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00617 107 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00616 534 107 108 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00615 105 104 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00614 534 105 106 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00613 534 102 96 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00612 96 102 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00611 99 101 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00610 534 96 82 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00609 82 79 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00608 534 488 79 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00607 83 82 92 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00606 534 133 83 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00605 87 134 90 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00604 534 86 87 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00603 74 73 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00602 534 204 73 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00601 73 182 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00600 81 91 84 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00599 534 82 81 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00598 136 84 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00597 534 136 69 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00596 68 162 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00595 69 118 68 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00594 76 96 77 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00593 534 488 76 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00592 86 77 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00591 534 62 58 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00590 61 57 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00589 61 60 62 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00588 62 205 61 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00587 534 66 60 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00586 65 112 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00585 65 72 66 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00584 66 201 65 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00583 534 136 72 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00582 71 162 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00581 72 74 71 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00580 534 192 59 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00579 57 59 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00578 534 201 59 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00577 59 69 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00576 6 134 30 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00575 534 488 6 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00574 8 91 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00573 37 42 8 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00572 38 43 37 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00571 36 43 9 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00570 9 38 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00569 10 42 36 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00568 43 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00567 534 43 42 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00566 41 39 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00565 534 41 10 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00564 534 37 91 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00563 91 37 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00562 38 36 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00561 89 91 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00560 7 89 31 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00559 7 29 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00558 534 91 7 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00557 31 30 7 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00556 39 31 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00555 22 23 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00554 534 205 23 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00553 5 86 29 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00552 534 133 5 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00551 25 24 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00550 534 204 24 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00549 4 89 26 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00548 534 86 4 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00547 27 28 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00546 534 182 28 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00545 162 26 534 534 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00544 20 21 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00543 534 201 21 534 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00542 1 201 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00541 11 18 1 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00540 13 19 11 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00539 14 19 3 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00538 3 13 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00537 2 18 14 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00536 19 515 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00535 534 19 18 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00534 17 58 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00533 534 17 2 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00532 534 11 201 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00531 201 11 534 534 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00530 13 14 534 534 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00529 487 526 525 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00528 526 528 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00527 529 528 485 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00526 487 529 527 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00525 485 532 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00524 487 520 521 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00523 520 519 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00522 487 533 530 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00521 533 531 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00520 487 531 532 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00519 487 490 493 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00518 487 491 492 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00517 491 489 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00516 462 516 510 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00515 487 508 462 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00514 510 518 511 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00513 487 511 468 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00512 468 518 513 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00511 513 516 467 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00510 518 516 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00509 487 515 516 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00508 467 517 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00507 487 514 517 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00506 508 510 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00505 487 510 508 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00504 511 513 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00503 487 505 506 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00502 505 504 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00501 487 523 524 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00500 523 522 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00499 500 499 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00498 487 508 500 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00497 487 502 503 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00496 502 508 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00495 487 497 514 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00494 487 495 453 487 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00493 453 500 487 487 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00492 497 494 452 487 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00491 452 493 487 487 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00490 453 504 497 487 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00489 487 488 494 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00488 487 486 479 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00487 479 477 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00486 479 478 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00485 486 528 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00484 487 532 486 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00483 482 484 483 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00482 483 527 482 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00481 487 480 483 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00480 481 482 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00479 487 528 484 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00478 484 522 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00477 484 532 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00476 487 531 475 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00475 475 474 478 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00474 478 476 473 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00473 473 522 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00472 487 522 474 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00471 476 531 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00470 455 454 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00469 455 504 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00468 487 499 455 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00467 487 455 457 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00466 458 456 469 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00465 469 459 458 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00464 458 457 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00463 460 470 461 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00462 487 504 460 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00461 461 472 463 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00460 487 463 466 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00459 466 472 464 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00458 464 470 465 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00457 472 470 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00456 487 515 470 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00455 465 471 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00454 487 469 471 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00453 504 461 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00452 487 461 504 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00451 463 464 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00450 454 508 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00449 487 447 454 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00448 490 450 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00447 450 504 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00446 487 451 450 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00445 495 451 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00444 487 456 495 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00443 487 490 449 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00442 449 446 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00441 448 456 449 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00440 449 447 448 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00439 487 489 447 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00438 487 504 459 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00437 378 427 419 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00436 487 522 378 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00435 419 426 420 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00434 487 420 383 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00433 383 426 422 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00432 422 427 387 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00431 426 427 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00430 487 515 427 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00429 387 424 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00428 487 423 424 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00427 522 419 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00426 487 419 522 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00425 420 422 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00424 411 477 372 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00423 487 411 412 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00422 372 522 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00421 487 417 423 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00420 487 479 376 487 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00419 376 412 487 487 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00418 417 413 375 487 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00417 375 522 487 487 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00416 376 414 417 487 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00415 353 451 352 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00414 487 396 351 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00413 352 459 397 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00412 351 489 353 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00411 487 397 409 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00410 413 488 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00409 487 409 413 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00408 408 494 366 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00407 487 408 414 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00406 366 409 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00405 487 508 451 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00404 400 390 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00403 487 448 390 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00402 342 389 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00401 390 504 342 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00400 392 451 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00399 392 489 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00398 487 499 392 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00397 487 392 393 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00396 356 405 398 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00395 487 489 356 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00394 398 406 401 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00393 487 401 360 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00392 360 406 402 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00391 402 405 361 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00390 406 405 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00389 487 515 405 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00388 361 407 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00387 487 400 407 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00386 489 398 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00385 487 398 489 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00384 401 402 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00383 487 494 336 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00382 336 489 446 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00381 341 508 389 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00380 389 446 341 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00379 341 393 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00378 370 477 374 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00377 487 370 371 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00376 374 528 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00375 331 386 377 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00374 487 528 331 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00373 377 380 382 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00372 487 382 381 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00371 381 380 379 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00370 379 386 334 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00369 380 386 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00368 487 515 386 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00367 334 384 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00366 487 385 384 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00365 528 377 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00364 487 377 528 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00363 382 379 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00362 322 365 362 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00361 487 414 322 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00360 321 413 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00359 362 531 321 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00358 487 362 363 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00357 317 354 345 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00356 487 531 317 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00355 345 348 350 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00354 487 350 349 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00353 349 348 347 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00352 347 354 319 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00351 348 354 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00350 487 515 354 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00349 319 355 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00348 487 363 355 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00347 531 345 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00346 487 345 531 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00345 350 347 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00344 487 373 385 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00343 487 481 328 487 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00342 328 371 487 487 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00341 373 413 327 487 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00340 327 528 487 487 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00339 328 414 373 487 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00338 344 477 456 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00337 456 343 344 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00336 344 494 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00335 367 396 368 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00334 487 367 369 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00333 368 494 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00332 357 480 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00331 487 531 358 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00330 359 358 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00329 365 357 359 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00328 364 531 365 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00327 487 480 364 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00326 487 346 396 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00325 487 335 337 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00324 335 340 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00323 312 488 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00322 487 337 312 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00321 325 488 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00320 487 396 325 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00319 487 338 343 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00318 338 346 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00317 487 339 313 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00316 313 340 346 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00315 249 292 285 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00314 487 519 249 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00313 285 289 286 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00312 487 286 248 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00311 248 289 291 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00310 291 292 250 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00309 289 292 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00308 487 515 292 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00307 250 290 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00306 487 297 290 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00305 519 285 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00304 487 285 519 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00303 286 291 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00302 487 296 297 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00301 487 300 253 487 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00300 253 304 487 487 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00299 296 325 256 487 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00298 256 519 487 487 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00297 253 369 296 487 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00296 487 519 262 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00295 262 306 309 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00294 309 308 261 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00293 261 307 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00292 487 307 306 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00291 308 519 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00290 305 519 260 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00289 487 305 304 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00288 260 303 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00287 487 369 293 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00286 294 293 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00285 487 299 294 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00284 487 282 278 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00283 278 488 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00282 278 277 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00281 487 283 477 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00280 283 281 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00279 487 278 243 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00278 243 274 499 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00277 301 309 255 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00276 487 301 300 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00275 255 299 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00274 487 339 282 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00273 239 273 264 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00272 487 339 239 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00271 264 270 265 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00270 487 265 238 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00269 238 270 269 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00268 269 273 241 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00267 270 273 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00266 487 515 273 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00265 241 267 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00264 487 272 267 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00263 339 264 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00262 487 264 339 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00261 265 269 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00260 272 275 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00259 487 271 275 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00258 242 339 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00257 275 312 242 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00256 487 480 281 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00255 228 235 257 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00254 487 307 228 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00253 257 234 258 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00252 487 258 231 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00251 231 234 259 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00250 259 235 236 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00249 234 235 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00248 487 515 235 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00247 236 233 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00246 487 232 233 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00245 307 257 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00244 487 257 307 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00243 258 259 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00242 487 325 227 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00241 227 307 252 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00240 487 307 254 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00239 252 254 226 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00238 226 294 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00237 232 252 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00236 221 307 251 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00235 487 294 221 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00234 222 325 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00233 251 299 222 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00232 487 251 220 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00231 214 219 245 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00230 487 299 214 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00229 245 216 246 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00228 487 246 213 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00227 213 216 247 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00226 247 219 218 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00225 216 219 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00224 487 515 219 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00223 218 217 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00222 487 220 217 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00221 299 245 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00220 487 245 299 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00219 246 247 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00218 487 488 197 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00217 197 339 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00216 197 277 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00215 487 240 271 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00214 200 197 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00213 199 202 200 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00212 240 210 199 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00211 274 281 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00210 487 206 274 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00209 487 204 274 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00208 274 205 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00207 487 244 210 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00206 244 211 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00205 487 205 192 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00204 487 237 340 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00203 193 203 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00202 194 192 193 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00201 237 201 194 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00200 487 201 206 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00199 202 205 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00198 487 206 202 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00197 487 191 480 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00196 480 303 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00195 480 307 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00194 170 182 153 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00193 487 170 203 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00192 153 211 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00191 487 184 185 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00190 184 299 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00189 487 299 303 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00188 487 186 187 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00187 186 307 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00186 487 519 191 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00185 487 182 277 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00184 487 169 204 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00183 169 171 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00182 165 210 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00181 165 162 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00180 487 205 165 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00179 487 165 167 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00178 487 168 152 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00177 152 166 151 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00176 151 167 177 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00175 155 183 175 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00174 487 171 155 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00173 175 178 173 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00172 487 173 154 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00171 154 178 180 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00170 180 183 156 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00169 178 183 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00168 487 515 183 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00167 156 179 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00166 487 177 179 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00165 171 175 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00164 487 175 171 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00163 173 180 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00162 487 201 150 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00161 150 210 157 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00160 160 192 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00159 160 158 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00158 487 204 160 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00157 487 160 166 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00156 487 171 211 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00155 211 171 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00154 487 119 118 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00153 119 203 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00152 138 144 140 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00151 487 182 138 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00150 140 147 139 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00149 487 139 142 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00148 142 147 141 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00147 141 144 146 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00146 147 144 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00145 487 515 144 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00144 146 145 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00143 487 143 145 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00142 182 140 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00141 487 140 182 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00140 139 141 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00139 487 148 149 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00138 148 339 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00137 487 133 134 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00136 113 162 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00135 487 277 113 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00134 135 132 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00133 132 162 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00132 487 182 132 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00131 487 135 131 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00130 131 136 130 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00129 137 136 143 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00128 143 277 137 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00127 137 135 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00126 487 130 117 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 117 204 168 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00124 120 129 124 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00123 487 205 120 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00122 124 128 121 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00121 487 121 123 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00120 123 128 122 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00119 122 129 127 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00118 128 129 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00117 487 515 129 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00116 127 126 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00115 487 125 126 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00114 205 124 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00113 487 124 205 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00112 121 122 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00111 487 110 114 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00110 111 113 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00109 109 157 111 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00108 110 192 109 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00107 487 113 158 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00106 487 158 112 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00105 112 201 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00104 112 210 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00103 125 115 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 487 114 115 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00101 116 205 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00100 115 130 116 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00099 53 89 93 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00098 487 92 53 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00097 52 90 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00096 93 91 52 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00095 487 93 104 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00094 54 107 102 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00093 487 96 54 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00092 102 108 99 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00091 487 99 55 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00090 55 108 101 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00089 101 107 56 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00088 108 107 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00087 487 515 107 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00086 56 105 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00085 487 104 105 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00084 96 102 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00083 487 102 96 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00082 99 101 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00081 79 488 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00080 51 96 82 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00079 487 79 51 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00078 92 133 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00077 487 82 92 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00076 90 86 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00075 487 134 90 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00074 73 182 50 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 487 73 74 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 50 204 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 136 84 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 84 82 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00069 487 91 84 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00068 48 162 69 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 69 118 48 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 48 136 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00065 86 77 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00064 77 488 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00063 487 96 77 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00062 58 62 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00061 487 57 62 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00060 46 60 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00059 62 205 46 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00058 60 66 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00057 487 112 66 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00056 47 72 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00055 66 201 47 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00054 49 162 72 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 72 74 49 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00052 49 136 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00051 487 59 57 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 45 192 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 44 69 45 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 59 201 44 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 30 488 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00046 487 134 30 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 34 43 37 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00044 487 91 34 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00043 37 42 38 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00042 487 38 35 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00041 35 42 36 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00040 36 43 40 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00039 42 43 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00038 487 515 43 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00037 40 41 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00036 487 39 41 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00035 91 37 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00034 487 37 91 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00033 38 36 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00032 487 91 89 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 32 89 31 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00030 487 30 32 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00029 33 29 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00028 31 91 33 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00027 487 31 39 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 487 23 22 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 23 205 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00024 29 133 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00023 487 86 29 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00022 487 24 25 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 24 204 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00020 26 86 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00019 487 89 26 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00018 487 28 27 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00017 28 182 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00016 487 26 162 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00015 487 21 20 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00014 21 201 487 487 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00013 12 19 11 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00012 487 201 12 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00011 11 18 13 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00010 487 13 16 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00009 16 18 14 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00008 14 19 15 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00007 18 19 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00006 487 515 19 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 15 17 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 487 58 17 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00003 201 11 487 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 487 11 201 487 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 13 14 487 487 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
C537 7 487 7.43e-15
C532 11 487 2.871e-14
C530 13 487 2.005e-14
C529 14 487 2.632e-14
C526 17 487 2.321e-14
C525 18 487 4.869e-14
C524 19 487 5.165e-14
C523 20 487 3.624e-14
C522 21 487 1.568e-14
C521 22 487 5.736e-14
C520 23 487 1.568e-14
C519 24 487 1.568e-14
C518 25 487 3.624e-14
C517 26 487 5.331e-14
C516 27 487 2.928e-14
C515 28 487 1.568e-14
C514 29 487 7.201e-14
C513 30 487 5.521e-14
C512 31 487 2.445e-14
C507 36 487 2.632e-14
C506 37 487 2.871e-14
C505 38 487 2.005e-14
C504 39 487 7.034e-14
C502 41 487 2.321e-14
C501 42 487 4.869e-14
C500 43 487 5.165e-14
C495 48 487 4.11e-15
C494 49 487 4.11e-15
C485 57 487 6.101e-14
C484 58 487 6.078e-14
C483 59 487 2.605e-14
C482 60 487 4.637e-14
C481 61 487 6.05e-15
C480 62 487 1.767e-14
C477 65 487 6.05e-15
C476 66 487 1.767e-14
C473 69 487 6.317e-14
C472 70 487 6.05e-15
C470 72 487 5.417e-14
C469 73 487 1.8635e-14
C468 74 487 4.633e-14
C465 77 487 1.8635e-14
C463 79 487 1.662e-14
C460 82 487 8.473e-14
C458 84 487 1.8635e-14
C456 86 487 1.4014e-13
C453 89 487 1.3676e-13
C452 90 487 5.041e-14
C451 91 487 1.7952e-13
C450 92 487 6.241e-14
C449 93 487 2.445e-14
C448 94 487 7.43e-15
C446 96 487 1.3565e-13
C443 99 487 2.005e-14
C441 101 487 2.632e-14
C440 102 487 2.871e-14
C438 104 487 7.034e-14
C437 105 487 2.321e-14
C435 107 487 5.165e-14
C434 108 487 4.869e-14
C431 110 487 2.605e-14
C429 112 487 6.213e-14
C428 113 487 8.482e-14
C427 114 487 7.661e-14
C426 115 487 1.767e-14
C423 118 487 5.713e-14
C422 119 487 1.568e-14
C420 121 487 2.005e-14
C419 122 487 2.632e-14
C417 124 487 2.871e-14
C416 125 487 7.998e-14
C415 126 487 2.321e-14
C413 128 487 4.869e-14
C412 129 487 5.165e-14
C411 130 487 1.0658e-13
C409 132 487 1.8635e-14
C408 133 487 1.8991e-13
C407 134 487 8.596e-14
C406 135 487 8.852e-14
C405 136 487 1.9275e-13
C404 137 487 4.11e-15
C402 139 487 2.005e-14
C401 140 487 2.871e-14
C400 141 487 2.632e-14
C398 143 487 6.378e-14
C397 144 487 5.165e-14
C396 145 487 2.321e-14
C394 147 487 4.869e-14
C393 148 487 1.568e-14
C392 149 487 5.328e-14
C383 157 487 4.863e-14
C382 158 487 7.645e-14
C380 160 487 2.455e-14
C378 162 487 2.347e-13
C375 165 487 2.455e-14
C374 166 487 7.152e-14
C373 167 487 5.852e-14
C372 168 487 5.513e-14
C371 169 487 1.568e-14
C370 170 487 1.8635e-14
C369 171 487 1.1828e-13
C367 173 487 2.005e-14
C365 175 487 2.871e-14
C363 177 487 9.226e-14
C362 178 487 4.869e-14
C361 179 487 2.321e-14
C360 180 487 2.632e-14
C358 182 487 2.5829e-13
C357 183 487 5.165e-14
C356 184 487 1.568e-14
C355 185 487 6.24e-14
C354 186 487 1.568e-14
C353 187 487 6.24e-14
C349 191 487 5.064e-14
C348 192 487 1.6034e-13
C343 197 487 5.047e-14
C339 201 487 3.1917e-13
C338 202 487 4.741e-14
C337 203 487 1.3132e-13
C336 204 487 2.3063e-13
C335 205 487 3.1753e-13
C334 206 487 7.48e-14
C330 210 487 1.8294e-13
C329 211 487 9.574e-14
C324 216 487 4.869e-14
C323 217 487 2.321e-14
C321 219 487 5.165e-14
C320 220 487 5.234e-14
C317 223 487 7.43e-15
C308 232 487 7.062e-14
C306 233 487 2.321e-14
C305 234 487 4.869e-14
C304 235 487 5.165e-14
C302 237 487 2.605e-14
C299 240 487 2.605e-14
C295 244 487 1.568e-14
C294 245 487 2.871e-14
C293 246 487 2.005e-14
C292 247 487 2.632e-14
C288 251 487 2.445e-14
C287 252 487 1.932e-14
C286 253 487 4.11e-15
C285 254 487 2.356e-14
C282 257 487 2.871e-14
C281 258 487 2.005e-14
C280 259 487 2.632e-14
C274 264 487 2.871e-14
C273 265 487 2.005e-14
C271 267 487 2.321e-14
C269 269 487 2.632e-14
C268 270 487 4.869e-14
C267 271 487 6.461e-14
C266 272 487 5.358e-14
C265 273 487 5.165e-14
C264 274 487 6.786e-14
C263 275 487 1.767e-14
C262 276 487 6.05e-15
C261 277 487 2.6331e-13
C260 278 487 5.937e-14
C257 281 487 9.497e-14
C256 282 487 4.824e-14
C255 283 487 1.568e-14
C253 285 487 2.871e-14
C252 286 487 2.005e-14
C249 289 487 4.869e-14
C248 290 487 2.321e-14
C247 291 487 2.632e-14
C246 292 487 5.165e-14
C245 293 487 1.677e-14
C244 294 487 9.363e-14
C242 296 487 2.299e-14
C241 297 487 6.13e-14
C239 299 487 2.5506e-13
C238 300 487 4.258e-14
C237 301 487 1.8635e-14
C236 302 487 8.58e-15
C235 303 487 1.0846e-13
C234 304 487 5.158e-14
C233 305 487 1.8635e-14
C232 306 487 2.596e-14
C231 307 487 2.3941e-13
C230 308 487 2.16e-14
C229 309 487 5.675e-14
C228 310 487 7.76e-15
C226 312 487 6.927e-14
C218 320 487 9.7e-15
C215 323 487 7.43e-15
C213 325 487 1.3247e-13
C210 328 487 4.11e-15
C209 329 487 8.58e-15
C202 335 487 1.568e-14
C200 337 487 4.798e-14
C199 338 487 1.568e-14
C198 339 487 3.4353e-13
C197 340 487 1.0883e-13
C196 341 487 4.11e-15
C194 343 487 4.873e-14
C193 344 487 4.11e-15
C192 345 487 2.871e-14
C191 346 487 8.786e-14
C190 347 487 2.632e-14
C189 348 487 4.869e-14
C187 350 487 2.005e-14
C183 354 487 5.165e-14
C182 355 487 2.321e-14
C180 357 487 2.16e-14
C179 358 487 2.596e-14
C175 362 487 2.445e-14
C174 363 487 6.074e-14
C172 365 487 5.485e-14
C170 367 487 1.8635e-14
C168 369 487 9.649e-14
C167 370 487 1.8635e-14
C166 371 487 4.438e-14
C164 373 487 2.299e-14
C161 376 487 4.11e-15
C160 377 487 2.871e-14
C158 379 487 2.632e-14
C157 380 487 4.869e-14
C155 382 487 2.005e-14
C153 384 487 2.321e-14
C152 385 487 6.85e-14
C151 386 487 5.165e-14
C147 389 487 4.937e-14
C146 390 487 1.767e-14
C145 391 487 6.05e-15
C144 392 487 2.455e-14
C143 393 487 6.227e-14
C140 396 487 1.5523e-13
C139 397 487 2.306e-14
C138 398 487 2.871e-14
C136 400 487 8.958e-14
C135 401 487 2.005e-14
C134 402 487 2.632e-14
C131 405 487 5.165e-14
C130 406 487 4.869e-14
C129 407 487 2.321e-14
C128 408 487 1.8635e-14
C127 409 487 1.2783e-13
C125 411 487 1.8635e-14
C124 412 487 4.678e-14
C123 413 487 1.3059e-13
C122 414 487 1.3185e-13
C121 415 487 8.58e-15
C119 417 487 2.299e-14
C117 419 487 2.871e-14
C116 420 487 2.005e-14
C114 422 487 2.632e-14
C113 423 487 7.21e-14
C112 424 487 2.321e-14
C110 426 487 4.869e-14
C109 427 487 5.165e-14
C97 439 487 7.76e-15
C89 446 487 8.275e-14
C88 447 487 7.345e-14
C87 448 487 5.533e-14
C86 449 487 7.43e-15
C85 450 487 1.8635e-14
C84 451 487 1.3208e-13
C82 453 487 4.11e-15
C81 454 487 7.411e-14
C80 455 487 2.455e-14
C79 456 487 1.3354e-13
C78 457 487 5.987e-14
C77 458 487 4.11e-15
C76 459 487 9.148e-14
C74 461 487 2.871e-14
C72 463 487 2.005e-14
C71 464 487 2.632e-14
C66 469 487 6.738e-14
C65 470 487 5.165e-14
C64 471 487 2.321e-14
C63 472 487 4.869e-14
C61 474 487 2.596e-14
C59 476 487 2.16e-14
C58 477 487 2.0774e-13
C57 478 487 5.274e-14
C56 479 487 5.362e-14
C55 480 487 2.5977e-13
C54 481 487 6.542e-14
C53 482 487 1.853e-14
C52 483 487 4.11e-15
C51 484 487 5.377e-14
C49 486 487 7.216e-14
C48 487 487 6.02665e-12
C47 488 487 4.9918e-13
C46 489 487 2.4521e-13
C45 490 487 8.177e-14
C44 491 487 1.568e-14
C43 492 487 4.248e-14
C42 493 487 5.604e-14
C41 494 487 2.9941e-13
C40 495 487 4.786e-14
C39 496 487 8.58e-15
C38 497 487 2.299e-14
C36 499 487 1.547e-13
C35 500 487 4.966e-14
C33 502 487 1.568e-14
C32 503 487 3.288e-14
C31 504 487 2.5983e-13
C30 505 487 1.568e-14
C29 506 487 3.168e-14
C27 508 487 2.5285e-13
C25 510 487 2.871e-14
C24 511 487 2.005e-14
C22 513 487 2.632e-14
C21 514 487 9.37e-14
C20 515 487 8.75439e-13
C19 516 487 5.165e-14
C18 517 487 2.321e-14
C17 518 487 4.869e-14
C16 519 487 3.0842e-13
C15 520 487 1.568e-14
C14 521 487 4.104e-14
C13 522 487 2.3798e-13
C12 523 487 1.568e-14
C11 524 487 3.168e-14
C10 525 487 3.048e-14
C9 526 487 1.568e-14
C8 527 487 5.201e-14
C7 528 487 2.7609e-13
C6 529 487 1.8635e-14
C5 530 487 3.048e-14
C4 531 487 3.0231e-13
C3 532 487 1.2185e-13
C2 533 487 1.568e-14
C1 534 487 6.32402e-12
.ends cronometro_cougar

